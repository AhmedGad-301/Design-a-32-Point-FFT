`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/24/2022 08:25:57 PM
// Design Name: 
// Module Name: DFT2_TB
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
`define bits 16
`define CLOCK100 100
`define CLOCK20 20

module DFT2_TB;
    // Inputs
    reg                 clk_100,clk_20,reset;
    reg  [3:0]          enable;
    reg  [1:0]          SEL;
    reg  [31:0]         in08,in18,in28,in38,in48,in58,in68,in78,in88,in98,in108,in118,in128,in138,
                        in148,in158,in168,in178,in188,in198,in208,in218,in228,in238,in248,in258,
                        in268,in278,in288,in298,in308,in318;
    wire [(2*16)-1:0]   out0,out1,out2,out3,out4,out5,out6,out7,out8,out9,out10,out11,out12,out13,
                        out14,out15,out16,out17,out18,out19,out20,out21,out22,out23,out24,out25,
                        out26,out27,out28,out29,out30,out31;
    
    DFT_2_point #(7, 16) D2P (
    .clk_100(clk_100),
    .clk_50(clk_50),
    .reset(reset),
    .in0(in08),.in1(in18),.in2(in28),.in3(in38),.in4(in48),.in5(in58),.in6(in68),.in7(in78),
    .in8(in88),.in9(in98),.in10(in108),.in11(in118),.in12(in128),.in13(in138),.in14(in148),
    .in15(in158),.in16(in168),.in17(in178),.in18(in188),.in19(in198),.in20(in208),.in21(in218),
    .in22(in228),.in23(in238),.in24(in248),.in25(in258),.in26(in268),.in27(in278),.in28(in288),
    .in29(in298),.in30(in308),.in31(in318),
    .out0(out0),.out1(out1),.out2(out2),.out3(out3),.out4(out4),.out5(out5),.out6(out6),.out7(out7),
    .out8(out8),.out9(out9),.out10(out10),.out11(out11),.out12(out12),.out13(out13),.out14(out14),
    .out15(out15),.out16(out16),.out17(out17),.out18(out18),.out19(out19),.out20(out20),.out21(out21),
    .out22(out22),.out23(out23),.out24(out24),.out25(out25),.out26(out26),.out27(out27),.out28(out28),
    .out29(out29),.out30(out30),.out31(out31)
    );
    
    initial
        begin
            clk_100 = 1;
            clk_50 = 1;
            reset = 0;
            SEL = 0;
            enable = 0;
            in08 = 32'b000000000_0000000__000000001_0000000;
            in18 = 32'b000000000_0000000__000000001_0000000;
            in28 = 32'b000000000_0000000__000000001_0000000;
            in38 = 32'b000000000_0000000__000000001_0000000;
            in48 = 32'b000000000_0000000__000000001_0000000;
            in58 = 32'b000000000_0000000__000000001_0000000;
            in68 = 32'b000000000_0000000__000000001_0000000;
            in78 = 32'b000000000_0000000__000000001_0000000;
            in88 = 32'b000000000_0000000__000000001_0000000;
            in98 = 32'b000000000_0000000__000000001_0000000;
            in108 = 32'b000000000_0000000__000000001_0000000;
            in118 = 32'b000000000_0000000__000000001_0000000;
            in128 = 32'b000000000_0000000__000000001_0000000;
            in138 = 32'b000000000_0000000__000000001_0000000;
            in148 = 32'b000000000_0000000__000000001_0000000;
            in158 = 32'b000000000_0000000__000000001_0000000;
            in168 = 32'b000000000_0000000__000000001_0000000;
            in178 = 32'b000000000_0000000__000000001_0000000;
            in188 = 32'b000000000_0000000__000000001_0000000;
            in198 = 32'b000000000_0000000__000000001_0000000;
            in208 = 32'b000000000_0000000__000000001_0000000;
            in218 = 32'b000000000_0000000__000000001_0000000;
            in228 = 32'b000000000_0000000__000000001_0000000;
            in238 = 32'b000000000_0000000__000000001_0000000;
            in248 = 32'b000000000_0000000__000000001_0000000;
            in258 = 32'b000000000_0000000__000000001_0000000;
            in268 = 32'b000000000_0000000__000000001_0000000;
            in278 = 32'b000000000_0000000__000000001_0000000;
            in288 = 32'b000000000_0000000__000000001_0000000;
            in298 = 32'b000000000_0000000__000000001_0000000;
            in308 = 32'b000000000_0000000__000000001_0000000;
            in318 = 32'b000000000_0000000__000000001_0000000;
        end
    
    always #(500/`CLOCK100) clk_100 = !clk_100;
    always #(500/`CLOCK20) clk_20 = !clk_20;
endmodule
