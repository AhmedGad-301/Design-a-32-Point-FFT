`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/24/2022 02:18:40 AM
// Design Name: 
// Module Name: TOP_TB
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
`define CLOCK1 100
`define CLOCK2 20

module TOP_TB;
    
    reg                 clk_100,clk_20,reset;
    reg [7:0]           in08,in18,in28,in38,in48,in58,in68,in78,in88,in98,in108,in118,in128,in138,
                        in148,in158,in168,in178,in188,in198,in208,in218,in228,in238,in248,in258,
                        in268,in278,in288,in298,in308,in318;
    wire [(2*16)-1:0]   out0,out1,out2,out3,out4,out5,out6,out7,out8,out9,out10,out11,out12,out13,
                        out14,out15,out16,out17,out18,out19,out20,out21,out22,out23,out24,out25,
                        out26,out27,out28,out29,out30,out31;
    TOP #(7, 16) TP (
    .clk_100(clk_100),
    .clk_20(clk_20),
    .reset(reset),
    .in08(in08),.in18(in18),.in28(in28),.in38(in38),.in48(in48),.in58(in58),.in68(in68),.in78(in78),
    .in88(in88),.in98(in98),.in108(in108),.in118(in118),.in128(in128),.in138(in138),.in148(in148),
    .in158(in158),.in168(in168),.in178(in178),.in188(in188),.in198(in198),.in208(in208),.in218(in218),
    .in228(in228),.in238(in238),.in248(in248),.in258(in258),.in268(in268),.in278(in278),.in288(in288),
    .in298(in298),.in308(in308),.in318(in318),
    .out0(out0),.out1(out1),.out2(out2),.out3(out3),.out4(out4),.out5(out5),.out6(out6),.out7(out7),
    .out8(out8),.out9(out9),.out10(out10),.out11(out11),.out12(out12),.out13(out13),.out14(out14),
    .out15(out15),.out16(out16),.out17(out17),.out18(out18),.out19(out19),.out20(out20),.out21(out21),
    .out22(out22),.out23(out23),.out24(out24),.out25(out25),.out26(out26),.out27(out27),.out28(out28),
    .out29(out29),.out30(out30),.out31(out31)
    );
    
    initial
        begin
            clk_100 = 1;
            clk_20 = 1;
            reset = 0;
            #100
//            in08 = 8'b00000001;
//            in18 = 8'b00000001;
//            in28 = 8'b00000010;
//            in38 = 8'b00000011;
//            in48 = 8'b00000010;
//            in58 = 8'b00000001;
//            in68 = 8'b00000001;
//            in78 = 8'b00000010;
//            in88 = 8'b00000011;
//            in98 = 8'b00000010;
//            in108 = 8'b00000001;
//            in118 = 8'b00000001;
//            in128 = 8'b00000010;
//            in138 = 8'b00000011;
//            in148 = 8'b00000010;
//            in158 = 8'b00000001;
//            in168 = 8'b00000001;
//            in178 = 8'b00000010;
//            in188 = 8'b00000011;
//            in198 = 8'b00000010;
//            in208 = 8'b00000001;
//            in218 = 8'b00000001;
//            in228 = 8'b00000010;
//            in238 = 8'b00000011;
//            in248 = 8'b00000010;
//            in258 = 8'b00000001;
//            in268 = 8'b00000001;
//            in278 = 8'b00000010;
//            in288 = 8'b00000011;
//            in298 = 8'b00000010;
//            in308 = 8'b00000001;
//            in318 = 8'b00000001;
//            #50
//            in08 = 8'b00000001;
//            in18 = 8'b00000001;
//            in28 = 8'b00000001;
//            in38 = 8'b00000001;
//            in48 = 8'b00000001;
//            in58 = 8'b00000001;
//            in68 = 8'b00000001;
//            in78 = 8'b00000001;
//            in88 = 8'b00000001;
//            in98 = 8'b00000001;
//            in108 = 8'b00000001;
//            in118 = 8'b00000001;
//            in128 = 8'b00000001;
//            in138 = 8'b00000001;
//            in148 = 8'b00000001;
//            in158 = 8'b00000001;
//            in168 = 8'b00000001;
//            in178 = 8'b00000001;
//            in188 = 8'b00000001;
//            in198 = 8'b00000001;
//            in208 = 8'b00000001;
//            in218 = 8'b00000001;
//            in228 = 8'b00000001;
//            in238 = 8'b00000001;
//            in248 = 8'b00000001;
//            in258 = 8'b00000001;
//            in268 = 8'b00000001;
//            in278 = 8'b00000001;
//            in288 = 8'b00000001;
//            in298 = 8'b00000001;
//            in308 = 8'b00000001;
//            in318 = 8'b00000001;
//            #50
//            reset = 0;
            in08 = 8'b00000000;
            in18 = 8'b00000000;
            in28 = 8'b00000000;
            in38 = 8'b00000000;
            in48 = 8'b00000000;
            in58 = 8'b00000000;
            in68 = 8'b00000000;
            in78 = 8'b00000000;
            in88 = 8'b00000000;
            in98 = 8'b00000000;
            in108 = 8'b00000000;
            in118 = 8'b00000000;
            in128 = 8'b00000000;
            in138 = 8'b00000000;
            in148 = 8'b00000000;
            in158 = 8'b00000000;
            in168 = 8'b00000000;
            in178 = 8'b00000000;
            in188 = 8'b00000000;
            in198 = 8'b00000000;
            in208 = 8'b00000000;
            in218 = 8'b00000000;
            in228 = 8'b00000000;
            in238 = 8'b00000000;
            in248 = 8'b00000000;
            in258 = 8'b00000000;
            in268 = 8'b00000000;
            in278 = 8'b00000000;
            in288 = 8'b00000000;
            in298 = 8'b00000000;
            in308 = 8'b00000000;
            in318 = 8'b00000000;
            #50
            in08 = 8'b00000001;
            in18 = 8'b00000001;
            in28 = 8'b00000010;
            in38 = 8'b00000011;
            in48 = 8'b00000010;
            in58 = 8'b00000001;
            in68 = 8'b00000001;
            in78 = 8'b00000010;
            in88 = 8'b00000011;
            in98 = 8'b00000010;
            in108 = 8'b00000001;
            in118 = 8'b00000001;
            in128 = 8'b00000010;
            in138 = 8'b00000011;
            in148 = 8'b00000010;
            in158 = 8'b00000001;
            in168 = 8'b00000001;
            in178 = 8'b00000010;
            in188 = 8'b00000011;
            in198 = 8'b00000010;
            in208 = 8'b00000001;
            in218 = 8'b00000001;
            in228 = 8'b00000010;
            in238 = 8'b00000011;
            in248 = 8'b00000010;
            in258 = 8'b00000001;
            in268 = 8'b00000001;
            in278 = 8'b00000010;
            in288 = 8'b00000011;
            in298 = 8'b00000010;
            in308 = 8'b00000001;
            in318 = 8'b00000001;
            #50
            in08 = 8'b00000000;
            in18 = 8'b00000000;
            in28 = 8'b00000000;
            in38 = 8'b00000000;
            in48 = 8'b00000000;
            in58 = 8'b00000000;
            in68 = 8'b00000000;
            in78 = 8'b00000000;
            in88 = 8'b00000000;
            in98 = 8'b00000000;
            in108 = 8'b00000000;
            in118 = 8'b00000000;
            in128 = 8'b00000000;
            in138 = 8'b00000000;
            in148 = 8'b00000000;
            in158 = 8'b00000000;
            in168 = 8'b00000000;
            in178 = 8'b00000000;
            in188 = 8'b00000000;
            in198 = 8'b00000000;
            in208 = 8'b00000000;
            in218 = 8'b00000000;
            in228 = 8'b00000000;
            in238 = 8'b00000000;
            in248 = 8'b00000000;
            in258 = 8'b00000000;
            in268 = 8'b00000000;
            in278 = 8'b00000000;
            in288 = 8'b00000000;
            in298 = 8'b00000000;
            in308 = 8'b00000000;
            in318 = 8'b00000000;
        end
    
    always #(500/`CLOCK1) clk_100 = !clk_100;
    always #(500/`CLOCK2) clk_20 = !clk_20;
    
    always @ (posedge clk_20)
        begin
            in08 = in08 + 1;
            in18 = in18 + 1;
            in28 = in28 + 1;
            in38 = in38 + 1;
            in48 = in48 + 1;
            in58 = in58 + 1;
            in68 = in68 + 1;
            in78 = in78 + 1;
            in88 = in88 + 1;
            in98 = in98 + 1;
            in108 = in108 + 1;
            in118 = in118 + 1;
            in128 = in128 + 1;
            in138 = in138 + 1;
            in148 = in148 + 1;
            in158 = in158 + 1;
            in168 = in168 + 1;
            in178 = in178 + 1;
            in188 = in188 + 1;
            in198 = in198 + 1;
            in208 = in208 + 1;
            in218 = in218 + 1;
            in228 = in228 + 1;
            in238 = in238 + 1;
            in248 = in248 + 1;
            in258 = in258 + 1;
            in268 = in268 + 1;
            in278 = in278 + 1;
            in288 = in288 + 1;
            in298 = in298 + 1;
            in308 = in308 + 1;
            in318 = in318 + 1;
        end
    
endmodule
